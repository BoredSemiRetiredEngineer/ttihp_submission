

// Testbench for Silly Project


module testbench;
    

    // Connections

    reg clk;
    reg rst_n;
    reg [7:0] ui_in;
   // reg [7:0] uio_in;
    wire [7:0] uo_out;

    silly1 silly1(.clk(clk), .rst_n(rst_n), .ui_in(ui_in), .uo_out(uo_out));

    initial 
        clk = 0;
     
    always
        #5 clk = ~clk;
    
    initial begin
        $dumpfile("tb_waveform.vcd");
        $dumpvars(0,testbench);
        #1 rst_n = 0;
        #2  ui_in = 8'h01;
        #10 ui_in = 8'h02;
        #20  ui_in = 8'h03;
        #30 ui_in = 8'h04;
        #40  ui_in = 8'h05;
        #50 ui_in = 8'h06;
        #60  ui_in = 8'h07;
        #70 ui_in = 8'h08;
        #80  ui_in = 8'h09;
        #90 ui_in = 8'h0A;
        #100  ui_in = 8'h0B;
        #110 ui_in = 8'h0C;
        #120  ui_in = 8'h0D;
        #130 ui_in = 8'h0E;
        #140  ui_in = 8'h0F;
        #150 ui_in = 8'h10;
        #160  ui_in = 8'h11;
        #170 ui_in = 8'h12;
        #180  ui_in = 8'h13;
        #190 ui_in = 8'h14;
        #200  ui_in = 8'h15;
        #210 ui_in = 8'h16;
        #220  ui_in = 8'h17;
        #230 ui_in = 8'h18;
        #240  ui_in = 8'h19;
        #250 ui_in = 8'h1A;
        #260  ui_in = 8'h1B;
        #270 ui_in = 8'h1C;
        #280  ui_in = 8'h1D;
        #290 ui_in = 8'h1E;
        #300  ui_in = 8'h1F;
        #310 ui_in = 8'h20;
        #320  ui_in = 8'h21;
        #320 ui_in = 8'h22;
        #340  ui_in = 8'h23;
        #350 ui_in = 8'h24;
        #360  ui_in = 8'h25;
        #370 ui_in = 8'h26;
        #380  ui_in = 8'h27;
        #390 ui_in = 8'h28;
        #400  ui_in = 8'h29;
        #410 ui_in = 8'h2A;
        #420  ui_in = 8'h2B;
        #430 ui_in = 8'h2C;
        #440  ui_in = 8'h2D;
        #450 ui_in = 8'h2E;
        #460  ui_in = 8'h2F;
        #470 ui_in = 8'h30;
        #480  ui_in = 8'h31;
        #490 ui_in = 8'h32;
        #500  ui_in = 8'h33;
        #510 ui_in = 8'h34;
        #520  ui_in = 8'h35;
        #530 ui_in = 8'h36;
        #540  ui_in = 8'h37;
        #550 ui_in = 8'h38;
        #560  ui_in = 8'h39;
        #570 ui_in = 8'h3A;
        #580  ui_in = 8'h3B;
        #590 ui_in = 8'h3C;
        #600  ui_in = 8'h3D;
        #610 ui_in = 8'h3E;
        #620  ui_in = 8'h3F;
        #630 ui_in = 8'h40;
        #640  ui_in = 8'h41;
        #650 ui_in = 8'h42;
        #660  ui_in = 8'h43;
        #670 ui_in = 8'h44;
        #680  ui_in = 8'h45;
        #690 ui_in = 8'h46;
        #700  ui_in = 8'h47;
        #710 ui_in = 8'h48;
        #720  ui_in = 8'h49;
        #730 ui_in = 8'h4A;
        #740  ui_in = 8'h4B;
        #750 ui_in = 8'h4C;
        #760  ui_in = 8'h4D;
        #770 ui_in = 8'h4E;
        #780  ui_in = 8'h4F;
        #790 ui_in = 8'h50;
        #800  ui_in = 8'h51;
        #810 ui_in = 8'h52;
        #820  ui_in = 8'h53;
        #830 ui_in = 8'h54;
        #840  ui_in = 8'h55;
        #850 ui_in = 8'h56;
        #860  ui_in = 8'h57;
        #870 ui_in = 8'h58;
        #880  ui_in = 8'h59;
        #890 ui_in = 8'h5A;
        #900  ui_in = 8'h5B;
        #910 ui_in = 8'h5C;
        #920  ui_in = 8'h5D;
        #930 ui_in = 8'h5E;
        #940  ui_in = 8'h5F;
        #950 ui_in = 8'h60;
        #960  ui_in = 8'h61;
        #970 ui_in = 8'h62;
        #980  ui_in = 8'h63;
        #990 ui_in = 8'h64;
        #10000  ui_in = 8'h65;
        #10010 ui_in = 8'h66;
        #10020  ui_in = 8'h67;
        #10030 ui_in = 8'h68;
        #10040  ui_in = 8'h69;
        #10050 ui_in = 8'h6A;
        #10060  ui_in = 8'h6B;
        #10070 ui_in = 8'h6C;
        #10080  ui_in = 8'h6D;
        #10090 ui_in = 8'h6E;
        #20000  ui_in = 8'h6F;
        #20010 ui_in = 8'h70;
        #20020  ui_in = 8'h71;
        #20030 ui_in = 8'h72;
        #20040  ui_in = 8'h73;
        #20050 ui_in = 8'h74;
        #20060  ui_in = 8'h75;
        #20070 ui_in = 8'h76;
        #20080  ui_in = 8'h77;
        #20090 ui_in = 8'h78;
        #30000  ui_in = 8'h79;
        #30010 ui_in = 8'h7A;
        #30020  ui_in = 8'h7B;
        #30030 ui_in = 8'h7C;
        #30040  ui_in = 8'h7D;
        #30050 ui_in = 8'h7E;
        #30060  ui_in = 8'h7F;
        #30070 ui_in = 8'h80;
        #30080  ui_in = 8'h81;
        #30090 ui_in = 8'h82;
        #30100  ui_in = 8'h83;
        #30110 ui_in = 8'h84;
        #30120  ui_in = 8'h85;
        #30130 ui_in = 8'h86;
        #30140  ui_in = 8'h87;
        #30150 ui_in = 8'h88;
        #30160  ui_in = 8'h89;
        #30170 ui_in = 8'h8A;
        #30180  ui_in = 8'h8B;
        #30190 ui_in = 8'h8C;
        #30200  ui_in = 8'h8D;
        #30210 ui_in = 8'h8E;
        #30220  ui_in = 8'h8F;
        #30230 ui_in = 8'h90;
        #30240  ui_in = 8'h91;
        #30250 ui_in = 8'h92;
        #30260  ui_in = 8'h93;
        #30270 ui_in = 8'h94;
        #30280  ui_in = 8'h95;
        #30290 ui_in = 8'h96;
        #30300  ui_in = 8'h97;
        #30310 ui_in = 8'h98;
        #30320  ui_in = 8'h99;
        #30330 ui_in = 8'h9A;
        #30340  ui_in = 8'h9B;
        #30350 ui_in = 8'h9C;
        #30360  ui_in = 8'h9D;
        #30370 ui_in = 8'h9E;
        #30380  ui_in = 8'h9F;
        #30390 ui_in = 8'hA0;
        #30400  ui_in = 8'hA1;
        #30410 ui_in = 8'hA2;
        #30420  ui_in = 8'hA3;
        #30430 ui_in = 8'hA4;
        #30440  ui_in = 8'hA5;
        #30450 ui_in = 8'hA6;
        #30460  ui_in = 8'hA7;
        #30470 ui_in = 8'hA8;
        #30480  ui_in = 8'hA9;
        #30490 ui_in = 8'hAA;
        #30500  ui_in = 8'hAB;
        #30510 ui_in = 8'hAC;
        #30520  ui_in = 8'hAD;
        #30530 ui_in = 8'hAE;
        #30540  ui_in = 8'hAF;
        #30550 ui_in = 8'hB0;
        #30560  ui_in = 8'hB1;
        #30570 ui_in = 8'hB2;
        #30580  ui_in = 8'hB3;
        #30590 ui_in = 8'hB4;
        #30600  ui_in = 8'hB5;
        #30610 ui_in = 8'hB6;
        #30620  ui_in = 8'hB7;
        #30630 ui_in = 8'hB8;
        #30640  ui_in = 8'hB9;
        #30650 ui_in = 8'hBA;
        #30660  ui_in = 8'hBB;
        #30670 ui_in = 8'hBC;
        #30680  ui_in = 8'hBD;
        #30690 ui_in = 8'hBE;
        #30700  ui_in = 8'hBF;
        #30710 ui_in = 8'hC0;
        #30720  ui_in = 8'hC1;
        #30730 ui_in = 8'hC2;
        #30740  ui_in = 8'hC3;
        #30750 ui_in = 8'hC4;
        #30760  ui_in = 8'hC5;
        #30770 ui_in = 8'hC6;
        #30780  ui_in = 8'hC7;
        #30790 ui_in = 8'hC8;
        #30800  ui_in = 8'hC9;
        #30810 ui_in = 8'hCA;
        #30820  ui_in = 8'hCB;
        #30830 ui_in = 8'hCC;
        #30840  ui_in = 8'hCD;
        #30850 ui_in = 8'hCE;
        #30860  ui_in = 8'hCF;
        #30870 ui_in = 8'hD0;
        #30880  ui_in = 8'hD1;
        #30890 ui_in = 8'hD2;
        #30900  ui_in = 8'hD3;
        #30910 ui_in = 8'hD4;
        #30920  ui_in = 8'hD5;
        #30930 ui_in = 8'hD6;
        #30940  ui_in = 8'hD7;
        #30950 ui_in = 8'hD8;
        #30960  ui_in = 8'hD9;
        #30970 ui_in = 8'hDA;
        #30980  ui_in = 8'hDB;
        #30990 ui_in = 8'hDC;
        #31000  ui_in = 8'hDD;
        #31010 ui_in = 8'hDE;
        #31020  ui_in = 8'hDF;
        #31030 ui_in = 8'hE0;
        #31040  ui_in = 8'hE1;
        #31050 ui_in = 8'hE2;
        #31060  ui_in = 8'hE3;
        #31070 ui_in = 8'hE4;
        #31080  ui_in = 8'hE5;
        #31090 ui_in = 8'hE6;
        #31100  ui_in = 8'hE7;
        #31110 ui_in = 8'hE8;
        #31120  ui_in = 8'hE9;
        #31130 ui_in = 8'hEA;
        #31140  ui_in = 8'hEB;
        #31150 ui_in = 8'hEC;
        #31160  ui_in = 8'hED;
        #31170 ui_in = 8'hEE;
        #31180  ui_in = 8'hEF;
        #31190 ui_in = 8'hF0;
        #31200  ui_in = 8'hF1;
        #31210 ui_in = 8'hF2;
        #31220  ui_in = 8'hF3;
        #31230 ui_in = 8'hF4;
        #31240  ui_in = 8'hF5;
        #31250 ui_in = 8'hF6;
        #31260  ui_in = 8'hF7;
        #31270 ui_in = 8'hF8;
        #31280  ui_in = 8'hF9;
        #31290 ui_in = 8'hFA;
        #31300  ui_in = 8'hFB;
        #31310 ui_in = 8'hFC;
        #31320  ui_in = 8'hFD;
        #31330 ui_in = 8'hFE;
        #31340  ui_in = 8'hFF;
        #40010 rst_n = ~rst_n;
        #40020 ui_in = 8'h01;
        #40030 ui_in = 8'h02;
        #40040  ui_in = 8'h03;
        #40050 ui_in = 8'h04;
        #40060  ui_in = 8'h05;
        #40070 ui_in = 8'h06;
        #40080  ui_in = 8'h07;
        #40090 ui_in = 8'h08;
        #40100  ui_in = 8'h09;
        #40110 ui_in = 8'h0A;
        #40120  ui_in = 8'h0B;
        #40130 ui_in = 8'h0C;
        #40140  ui_in = 8'h0D;
        #40150 ui_in = 8'h0E;
        #40160  ui_in = 8'h0F;
        #40170 ui_in = 8'h10;
        #40180  ui_in = 8'h11;
        #40190 ui_in = 8'h12;
        #40200  ui_in = 8'h13;
        #40210 ui_in = 8'h14;
        #40220  ui_in = 8'h15;
        #40230 ui_in = 8'h16;
        #40240  ui_in = 8'h17;
        #40250 ui_in = 8'h18;
        #40260  ui_in = 8'h19;
        #40270 ui_in = 8'h1A;
        #40280  ui_in = 8'h1B;
        #40290 ui_in = 8'h1C;
        #40300  ui_in = 8'h1D;
        #40310 ui_in = 8'h1E;
        #40320  ui_in = 8'h1F;
        #40330 ui_in = 8'h20;
        #40340  ui_in = 8'h21;
        #40350 ui_in = 8'h22;
        #40360  ui_in = 8'h23;
        #40370 ui_in = 8'h24;
        #40380  ui_in = 8'h25;
        #40390 ui_in = 8'h26;
        #40400  ui_in = 8'h27;
        #40410 ui_in = 8'h28;
        #40420  ui_in = 8'h29;
        #40430 ui_in = 8'h2A;
        #40440  ui_in = 8'h2B;
        #40450 ui_in = 8'h2C;
        #40460  ui_in = 8'h2D;
        #40470 ui_in = 8'h2E;
        #40480  ui_in = 8'h2F;
        #40490 ui_in = 8'h30;
        #40500  ui_in = 8'h31;
        #40510 ui_in = 8'h32;
        #40520  ui_in = 8'h33;
        #40530 ui_in = 8'h34;
        #40540  ui_in = 8'h35;
        #40550 ui_in = 8'h36;
        #40560  ui_in = 8'h37;
        #40570 ui_in = 8'h38;
        #40580  ui_in = 8'h39;
        #40590 ui_in = 8'h3A;
        #40600  ui_in = 8'h3B;
        #40610 ui_in = 8'h3C;
        #40620  ui_in = 8'h3D;
        #40630 ui_in = 8'h3E;
        #40640  ui_in = 8'h3F;
        #40650 ui_in = 8'h40;
        #40660  ui_in = 8'h41;
        #40670 ui_in = 8'h42;
        #40680  ui_in = 8'h43;
        #40690 ui_in = 8'h44;
        #40700  ui_in = 8'h45;
        #40710 ui_in = 8'h46;
        #40720  ui_in = 8'h47;
        #40730 ui_in = 8'h48;
        #40740  ui_in = 8'h49;
        #40750 ui_in = 8'h4A;
        #40760  ui_in = 8'h4B;
        #40770 ui_in = 8'h4C;
        #40780  ui_in = 8'h4D;
        #40790 ui_in = 8'h4E;
        #40800  ui_in = 8'h4F;
        #40810 ui_in = 8'h50;
        #40820  ui_in = 8'h51;
        #40830 ui_in = 8'h52;
        #40840  ui_in = 8'h53;
        #40850 ui_in = 8'h54;
        #40860  ui_in = 8'h55;
        #40870 ui_in = 8'h56;
        #40880  ui_in = 8'h57;
        #40890 ui_in = 8'h58;
        #40900  ui_in = 8'h59;
        #40910 ui_in = 8'h5A;
        #40920  ui_in = 8'h5B;
        #40930 ui_in = 8'h5C;
        #40940  ui_in = 8'h5D;
        #40950 ui_in = 8'h5E;
        #40960  ui_in = 8'h5F;
        #40970 ui_in = 8'h60;
        #40980  ui_in = 8'h61;
        #40990 ui_in = 8'h62;
        #41000  ui_in = 8'h63;
        #41010 ui_in = 8'h64;
        #41020  ui_in = 8'h65;
        #41030 ui_in = 8'h66;
        #41040  ui_in = 8'h67;
        #41050 ui_in = 8'h68;
        #41060  ui_in = 8'h69;
        #41070 ui_in = 8'h6A;
        #41080  ui_in = 8'h6B;
        #41090 ui_in = 8'h6C;
        #41000  ui_in = 8'h6D;
        #41010 ui_in = 8'h6E;
        #41020  ui_in = 8'h6F;
        #41030 ui_in = 8'h70;
        #41040  ui_in = 8'h71;
        #41050 ui_in = 8'h72;
        #41060  ui_in = 8'h73;
        #41070 ui_in = 8'h74;
        #41080  ui_in = 8'h75;
        #41090 ui_in = 8'h76;
        #41100  ui_in = 8'h77;
        #41110 ui_in = 8'h78;
        #41120  ui_in = 8'h79;
        #41130 ui_in = 8'h7A;
        #41140  ui_in = 8'h7B;
        #41150 ui_in = 8'h7C;
        #41160  ui_in = 8'h7D;
        #41170 ui_in = 8'h7E;
        #41180  ui_in = 8'h7F;
        #41190 ui_in = 8'h80;
        #41200  ui_in = 8'h81;
        #41210 ui_in = 8'h82;
        #41220  ui_in = 8'h83;
        #41230 ui_in = 8'h84;
        #41240  ui_in = 8'h85;
        #41250 ui_in = 8'h86;
        #41260  ui_in = 8'h87;
        #41270 ui_in = 8'h88;
        #41280  ui_in = 8'h89;
        #41290 ui_in = 8'h8A;
        #41300  ui_in = 8'h8B;
        #41310 ui_in = 8'h8C;
        #41320  ui_in = 8'h8D;
        #41330 ui_in = 8'h8E;
        #41340  ui_in = 8'h8F;
        #41350 ui_in = 8'h90;
        #41360  ui_in = 8'h91;
        #41370 ui_in = 8'h92;
        #41380  ui_in = 8'h93;
        #41390 ui_in = 8'h94;
        #41400  ui_in = 8'h95;
        #41410 ui_in = 8'h96;
        #41420  ui_in = 8'h97;
        #41430 ui_in = 8'h98;
        #41440  ui_in = 8'h99;
        #41450 ui_in = 8'h9A;
        #41460  ui_in = 8'h9B;
        #41470 ui_in = 8'h9C;
        #41480  ui_in = 8'h9D;
        #41490 ui_in = 8'h9E;
        #41500  ui_in = 8'h9F;
        #41510 ui_in = 8'hA0;
        #41520  ui_in = 8'hA1;
        #41530 ui_in = 8'hA2;
        #41540  ui_in = 8'hA3;
        #41550 ui_in = 8'hA4;
        #41560  ui_in = 8'hA5;
        #41570 ui_in = 8'hA6;
        #41580  ui_in = 8'hA7;
        #41590 ui_in = 8'hA8;
        #41600  ui_in = 8'hA9;
        #41610 ui_in = 8'hAA;
        #41620  ui_in = 8'hAB;
        #41630 ui_in = 8'hAC;
        #41640  ui_in = 8'hAD;
        #41650 ui_in = 8'hAE;
        #41660  ui_in = 8'hAF;
        #41670 ui_in = 8'hB0;
        #41680  ui_in = 8'hB1;
        #41690 ui_in = 8'hB2;
        #41700  ui_in = 8'hB3;
        #41710 ui_in = 8'hB4;
        #41720  ui_in = 8'hB5;
        #41730 ui_in = 8'hB6;
        #41740  ui_in = 8'hB7;
        #41750 ui_in = 8'hB8;
        #41760  ui_in = 8'hB9;
        #41770 ui_in = 8'hBA;
        #41780  ui_in = 8'hBB;
        #41790 ui_in = 8'hBC;
        #41800  ui_in = 8'hBD;
        #41810 ui_in = 8'hBE;
        #41820  ui_in = 8'hBF;
        #41830 ui_in = 8'hC0;
        #41840  ui_in = 8'hC1;
        #41850 ui_in = 8'hC2;
        #41860  ui_in = 8'hC3;
        #41870 ui_in = 8'hC4;
        #41880  ui_in = 8'hC5;
        #41890 ui_in = 8'hC6;
        #41900  ui_in = 8'hC7;
        #41910 ui_in = 8'hC8;
        #41920  ui_in = 8'hC9;
        #41930 ui_in = 8'hCA;
        #41940  ui_in = 8'hCB;
        #41950 ui_in = 8'hCC;
        #41960  ui_in = 8'hCD;
        #41970 ui_in = 8'hCE;
        #41980  ui_in = 8'hCF;
        #41990 ui_in = 8'hD0;
        #42000  ui_in = 8'hD1;
        #42010 ui_in = 8'hD2;
        #42020  ui_in = 8'hD3;
        #42030 ui_in = 8'hD4;
        #42040  ui_in = 8'hD5;
        #42050 ui_in = 8'hD6;
        #42060  ui_in = 8'hD7;
        #42070 ui_in = 8'hD8;
        #42080  ui_in = 8'hD9;
        #42090 ui_in = 8'hDA;
        #42100  ui_in = 8'hDB;
        #42110 ui_in = 8'hDC;
        #42120  ui_in = 8'hDD;
        #42130 ui_in = 8'hDE;
        #42140  ui_in = 8'hDF;
        #42150 ui_in = 8'hE0;
        #42160  ui_in = 8'hE1;
        #42170 ui_in = 8'hE2;
        #42180  ui_in = 8'hE3;
        #42190 ui_in = 8'hE4;
        #42200  ui_in = 8'hE5;
        #42210 ui_in = 8'hE6;
        #42220  ui_in = 8'hE7;
        #42230 ui_in = 8'hE8;
        #42240  ui_in = 8'hE9;
        #42250 ui_in = 8'hEA;
        #42260  ui_in = 8'hEB;
        #42270 ui_in = 8'hEC;
        #42280  ui_in = 8'hED;
        #42290 ui_in = 8'hEE;
        #42300  ui_in = 8'hEF;
        #42310 ui_in = 8'hF0;
        #42320  ui_in = 8'hF1;
        #42330 ui_in = 8'hF2;
        #42340  ui_in = 8'hF3;
        #42350 ui_in = 8'hF4;
        #42360  ui_in = 8'hF5;
        #42370 ui_in = 8'hF6;
        #42380  ui_in = 8'hF7;
        #42390 ui_in = 8'hF8;
        #42400  ui_in = 8'hF9;
        #42410 ui_in = 8'hFA;
        #42420  ui_in = 8'hFB;
        #42430 ui_in = 8'hFC;
        #42440  ui_in = 8'hFD;
        #42450 ui_in = 8'hFE;
        #42460  ui_in = 8'hFF;
        #45000 $finish;


    end
    initial begin
    $monitor("clk = %b, rst_n = %b : ui_in = %h, ==> uo_out = %h  ", clk, rst_n, ui_in, uo_out);
    end

endmodule
